module IF_ID(
    input wire clk,
    input wire rst,
    input wire[31:0] fe_pc,
    input wire[31:0] fe_inst,
    output reg[31:0] id_pc,
    output reg[31:0] id_inst
);

endmodule