`include "../defines.sv"
module decode(
);

endmodule