`include "../defines.sv"
module icache(
    input PC pc,
    output INST[1:0] inst
);

endmodule