`include "../defines.svh"
module decoder(
);

endmodule