`include "../includes/defines.v"
module IF(
    input wire rst,

    input wire[31:0] pc,
    input wire[31:0] pc_4,

    input wire[31:0] inst_1,
    input wire[31:0] inst_2
);



endmodule