`include "../defines.svh"
module issue(
    input ISSUE_QUEUE_ELEMENT [1:0] issue_require,
    input IQ_ADDR iq_size
);

score_board score_board0(

);

always_comb begin

end

endmodule