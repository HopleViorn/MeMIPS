`include "defines.sv"
module icache(
    input PC pc,
    output INST[3:0] inst
);

endmodule