module FIFO(
    input wire clk,
    input wire rst,
    input wire[31:0] inst1,
    input wire[31:0] inst2
);

endmodule