module IF(
    input wire clk,
    input wire rst,
    input wire[31:0] brunch_addr,
    input wire brucnflag,
    output reg[31:0] pc
);


endmodule