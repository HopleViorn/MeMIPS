`include "../defines.svh"
module decode(
);

endmodule