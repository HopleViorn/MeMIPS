module MeMIPS(

);


endmodule