module mips(
    input wire clk,
    input wire rst
);


endmodule