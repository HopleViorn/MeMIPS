`include "defines.svh"
module pc_select(

    output logic[31:0] pc
);

always_comb begin
    
end

endmodule