`include "../defines.svh"
module issue(
    
);

endmodule