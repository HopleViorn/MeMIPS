module ID(
    input wire rst,
    input wire[31:0] pc,
    input wire[31:0] inst
);

endmodule