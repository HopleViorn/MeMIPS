module pc_predictor(

);

endmodule