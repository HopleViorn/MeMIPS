module control(
);

endmodule