`include "../defines.svh"
module decoder(
    input INST inst
);

endmodule