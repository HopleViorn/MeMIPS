`include "../defines.svh"
module pc_select(
    input PC_CHECK pc_fetch,
    input PC_CHECK pc_execute,
    output logic[31:0] pc
);

always_comb begin
    
end

endmodule