module ID_EX(
    input wire clk,
    input wire rst
);

endmodule