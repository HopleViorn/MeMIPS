module IF(
    input wire clk,
    input wire rst,
    output reg[31:0] pc
);


endmodule