`include "../defines.sv"
module decoder(
    input INST inst
);

endmodule