module IF(
    input wire clk,
    input wire rst,
    input wire[31:0] brunch_addr,
    input wire brucn_flag,
    output reg[31:0] pc
);


endmodule