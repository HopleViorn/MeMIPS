module MeMIPS(

);
