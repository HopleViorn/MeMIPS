`include "../defines.sv"
module commmit(
    input CMT_REQUIRE cmt_require[1:0]
);

endmodule